// hazard unit

module hazard_unit (

);

endmodule